

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO top 
  PIN ROM_address[11] 
    ANTENNAPARTIALMETALAREA 8.2004 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 33.8604 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 65.2232 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 270.535 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 277.676 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1150.7 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 9.6712 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 40.3912 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 1.5337 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 462.048 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 1544.96 LAYER metal6 ;
  END ROM_address[11]
  PIN ROM_address[10] 
    ANTENNAPARTIALMETALAREA 0.6356 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6332 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 49.0784 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 203.65 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 291.334 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1207.28 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 9.4472 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 39.788 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 1.5337 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 383.04 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 1281.6 LAYER metal6 ;
  END ROM_address[10]
  PIN ROM_address[9] 
    ANTENNAPARTIALMETALAREA 0.728 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.016 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 24.3264 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 101.106 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 292.936 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1213.92 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 11.928 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 49.7408 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 1.5337 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 424.608 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 1420.16 LAYER metal6 ;
  END ROM_address[9]
  PIN ROM_address[8] 
    ANTENNAPARTIALMETALAREA 268.262 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1111.37 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 6.1824 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 25.9376 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 10.976 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 45.7968 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 10.8528 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 45.2864 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 1.5337 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 479.136 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 1601.92 LAYER metal6 ;
  END ROM_address[8]
  PIN ROM_address[7] 
    ANTENNAPARTIALMETALAREA 268.582 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1112.7 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.4368 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1344 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1368 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 1.5337 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 561.792 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 1877.44 LAYER metal6 ;
  END ROM_address[7]
  PIN ROM_address[6] 
    ANTENNAPARTIALMETALAREA 263.29 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1090.77 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 2.7272 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.6232 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNADIFFAREA 1.5337 LAYER metal4 ; 
    ANTENNAPARTIALMETALAREA 147.885 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 612.99 LAYER metal4 ;
  END ROM_address[6]
  PIN ROM_address[5] 
    ANTENNAPARTIALMETALAREA 264.79 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1096.99 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 3.7688 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.9384 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 116.76 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 484.045 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.5337 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 21.1288 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 87.8584 LAYER metal5 ;
  END ROM_address[5]
  PIN ROM_address[4] 
    ANTENNAPARTIALMETALAREA 266.067 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1102.28 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 2.9008 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.3424 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 123.973 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 513.926 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.5337 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 27.188 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 112.961 LAYER metal5 ;
  END ROM_address[4]
  PIN ROM_address[3] 
    ANTENNAPARTIALMETALAREA 273.33 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1132.37 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 18.9952 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 79.0192 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 99.8256 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 413.888 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.5337 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 30.8504 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 128.134 LAYER metal5 ;
  END ROM_address[3]
  PIN ROM_address[2] 
    ANTENNAPARTIALMETALAREA 412.359 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1708.34 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNADIFFAREA 1.5337 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 62.7424 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 260.258 LAYER metal3 ;
  END ROM_address[2]
  PIN ROM_address[1] 
    ANTENNADIFFAREA 1.5386 LAYER metal2 ; 
    ANTENNAPARTIALMETALAREA 149.064 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 618.199 LAYER metal2 ;
  END ROM_address[1]
  PIN ROM_address[0] 
    ANTENNADIFFAREA 1.5386 LAYER metal2 ; 
    ANTENNAPARTIALMETALAREA 148.747 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 616.888 LAYER metal2 ;
  END ROM_address[0]
  PIN ROM_out[31] 
    ANTENNAPARTIALMETALAREA 74.6592 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 309.627 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.5936 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1088 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal3 ; 
    ANTENNAMAXAREACAR 331.518 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 1370.51 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.500639 LAYER via3 ;
  END ROM_out[31]
  PIN ROM_out[30] 
    ANTENNAPARTIALMETALAREA 66.178 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 274.491 LAYER metal2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3618 LAYER metal2 ; 
    ANTENNAMAXAREACAR 184.66 LAYER metal2 ;
    ANTENNAMAXSIDEAREACAR 761.122 LAYER metal2 ;
    ANTENNAMAXCUTCAR 0.216694 LAYER via2 ;
  END ROM_out[30]
  PIN ROM_out[29] 
    ANTENNAPARTIALMETALAREA 7.5824 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 31.4128 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 22.344 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 92.8928 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.4368 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1344 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1704.29 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5685.76 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5458.08 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18220.4 LAYER metal6 ;
  END ROM_out[29]
  PIN ROM_out[28] 
    ANTENNAPARTIALMETALAREA 8.248 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 34.0576 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 24.2536 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 100.804 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4848 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1699.58 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5670.08 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5438.12 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18149.9 LAYER metal6 ;
  END ROM_out[28]
  PIN ROM_out[27] 
    ANTENNAPARTIALMETALAREA 0.3388 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4036 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 64.5288 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 267.658 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.5936 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.784 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.9912 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 4.4312 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1723.1 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5748.48 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5528.52 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18466.8 LAYER metal6 ;
  END ROM_out[27]
  PIN ROM_out[26] 
    ANTENNAPARTIALMETALAREA 0.8848 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.6656 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 28.1652 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 117.009 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.7504 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4336 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1731.17 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5775.36 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5537.02 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18478 LAYER metal6 ;
  END ROM_out[26]
  PIN ROM_out[25] 
    ANTENNAPARTIALMETALAREA 0.8924 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.5844 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 15.0528 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 62.6864 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.4368 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1344 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1749.07 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5844.64 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5611.02 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18771 LAYER metal6 ;
  END ROM_out[25]
  PIN ROM_out[24] 
    ANTENNAPARTIALMETALAREA 0.3528 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4616 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 28.2464 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 117.346 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.9072 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.0832 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1753.78 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5860.32 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5629.91 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18835 LAYER metal6 ;
  END ROM_out[24]
  PIN ROM_out[23] 
    ANTENNAPARTIALMETALAREA 0.9596 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.8628 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 9.324 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 38.9528 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.4368 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1344 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1743.79 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5827.04 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5599.69 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18735.7 LAYER metal6 ;
  END ROM_out[23]
  PIN ROM_out[22] 
    ANTENNAPARTIALMETALAREA 8.5652 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 35.4844 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 29.4448 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 122.31 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4848 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1368 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1703.62 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5683.52 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5449.33 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18185.9 LAYER metal6 ;
  END ROM_out[22]
  PIN ROM_out[21] 
    ANTENNAPARTIALMETALAREA 7.504 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 31.088 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 2.7272 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.6232 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4848 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1368 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1702.94 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5681.28 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5530.67 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18524.6 LAYER metal6 ;
  END ROM_out[21]
  PIN ROM_out[20] 
    ANTENNAPARTIALMETALAREA 2.9232 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.1104 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 5.4824 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 23.0376 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1368 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 1.512 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 6.5888 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1728.48 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5766.4 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5542.58 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18508 LAYER metal6 ;
  END ROM_out[20]
  PIN ROM_out[19] 
    ANTENNAPARTIALMETALAREA 0.728 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.016 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.392 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9488 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1368 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.9912 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 4.4312 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1733.18 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5782.08 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5541.97 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18493.3 LAYER metal6 ;
  END ROM_out[19]
  PIN ROM_out[18] 
    ANTENNAPARTIALMETALAREA 4.4688 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 18.5136 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 2.9008 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.3424 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4848 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1719.74 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5737.28 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5498.74 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18348.9 LAYER metal6 ;
  END ROM_out[18]
  PIN ROM_out[17] 
    ANTENNAPARTIALMETALAREA 4.3344 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.9568 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 8.6464 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 36.1456 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4848 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1736.4 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5802.4 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5563.04 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18602.9 LAYER metal6 ;
  END ROM_out[17]
  PIN ROM_out[16] 
    ANTENNAPARTIALMETALAREA 4.3344 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.9568 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 6.6192 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 27.7472 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4848 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1709.66 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5703.68 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5491.58 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18346.4 LAYER metal6 ;
  END ROM_out[16]
  PIN ROM_out[15] 
    ANTENNAPARTIALMETALAREA 0.4144 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7168 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 23.6544 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 98.3216 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.5936 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.784 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1735.87 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5791.04 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5549.01 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18515.5 LAYER metal6 ;
  END ROM_out[15]
  PIN ROM_out[14] 
    ANTENNAPARTIALMETALAREA 0.3444 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4268 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 25.9896 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 107.996 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.9072 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.0832 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1733.18 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5782.08 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5544.51 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18503.8 LAYER metal6 ;
  END ROM_out[14]
  PIN ROM_out[13] 
    ANTENNAPARTIALMETALAREA 7.5376 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 31.2272 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 33.9752 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 141.079 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4848 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1368 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1704.96 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5688 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5455.56 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18208.2 LAYER metal6 ;
  END ROM_out[13]
  PIN ROM_out[12] 
    ANTENNAPARTIALMETALAREA 7.784 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 32.248 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 22.12 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 91.9648 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4848 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1698.91 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5667.84 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5442.11 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18170.2 LAYER metal6 ;
  END ROM_out[12]
  PIN ROM_out[11] 
    ANTENNAPARTIALMETALAREA 7.9464 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 32.9208 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 13.3168 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 55.4944 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4848 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1368 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1700.26 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5672.32 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5452.91 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18210.5 LAYER metal6 ;
  END ROM_out[11]
  PIN ROM_out[10] 
    ANTENNAPARTIALMETALAREA 8.2508 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 34.0692 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 13.8376 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 57.652 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4848 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1368 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1703.62 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5683.52 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5460.53 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18233.3 LAYER metal6 ;
  END ROM_out[10]
  PIN ROM_out[9] 
    ANTENNAPARTIALMETALAREA 4.3344 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.9568 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 14.0168 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 58.7192 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 390.085 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1616.39 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 4.7096 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 20.4856 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal5 ; 
    ANTENNAMAXAREACAR 24.09 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 99.9923 LAYER metal5 ;
    ANTENNAMAXCUTCAR 1.00128 LAYER via5 ;
  END ROM_out[9]
  PIN ROM_out[8] 
    ANTENNAPARTIALMETALAREA 2.7664 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.4608 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 1.1872 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.2176 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal3 ; 
    ANTENNAMAXAREACAR 16.7414 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 69.5479 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.500639 LAYER via3 ;
  END ROM_out[8]
  PIN ROM_out[7] 
    ANTENNAPARTIALMETALAREA 146.308 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 606.46 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4848 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 4.6368 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 19.5344 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal5 ; 
    ANTENNAMAXAREACAR 26.4681 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 109.844 LAYER metal5 ;
    ANTENNAMAXCUTCAR 1.00128 LAYER via5 ;
  END ROM_out[7]
  PIN ROM_out[6] 
    ANTENNAPARTIALMETALAREA 5.572 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 24.708 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal3 ; 
    ANTENNAMAXAREACAR 28.4527 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 118.066 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.500639 LAYER via3 ;
  END ROM_out[6]
  PIN ROM_out[5] 
    ANTENNAPARTIALMETALAREA 1.2908 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.9972 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal3 ; 
    ANTENNAMAXAREACAR 13.675 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 53.7331 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.500639 LAYER via3 ;
  END ROM_out[5]
  PIN ROM_out[4] 
    ANTENNAPARTIALMETALAREA 1.9264 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.3056 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 4.5136 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 19.024 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal4 ; 
    ANTENNAMAXAREACAR 25.3059 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 103.992 LAYER metal4 ;
    ANTENNAMAXCUTCAR 0.750958 LAYER via4 ;
  END ROM_out[4]
  PIN ROM_out[3] 
    ANTENNAPARTIALMETALAREA 3.7324 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.762 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal3 ; 
    ANTENNAMAXAREACAR 16.9649 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 69.4368 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.500639 LAYER via3 ;
  END ROM_out[3]
  PIN ROM_out[2] 
    ANTENNAPARTIALMETALAREA 1.7472 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.5376 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal3 ; 
    ANTENNAMAXAREACAR 9.12452 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 36.9553 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.500639 LAYER via3 ;
  END ROM_out[2]
  PIN ROM_out[1] 
    ANTENNAPARTIALMETALAREA 1.9124 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.5724 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal3 ; 
    ANTENNAMAXAREACAR 15.159 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 60.9183 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.500639 LAYER via3 ;
  END ROM_out[1]
  PIN ROM_out[0] 
    ANTENNAPARTIALMETALAREA 174.255 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 722.239 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.56 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9696 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal4 ; 
    ANTENNAMAXAREACAR 16.2586 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 68.5849 LAYER metal4 ;
    ANTENNAMAXCUTCAR 0.750958 LAYER via4 ;
  END ROM_out[0]
  PIN DRAM_WEn[3] 
    ANTENNAPARTIALMETALAREA 199.976 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 828.472 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNADIFFAREA 3.6652 LAYER metal4 ; 
    ANTENNAPARTIALMETALAREA 215.723 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 894.035 LAYER metal4 ;
  END DRAM_WEn[3]
  PIN DRAM_WEn[2] 
    ANTENNAPARTIALMETALAREA 205.159 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 849.944 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNADIFFAREA 9.072 LAYER metal4 ; 
    ANTENNAPARTIALMETALAREA 193.178 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 800.632 LAYER metal4 ;
  END DRAM_WEn[2]
  PIN DRAM_WEn[1] 
    ANTENNAPARTIALMETALAREA 198.727 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 823.298 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNADIFFAREA 5.20755 LAYER metal4 ; 
    ANTENNAPARTIALMETALAREA 171.819 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 712.147 LAYER metal4 ;
  END DRAM_WEn[1]
  PIN DRAM_WEn[0] 
    ANTENNAPARTIALMETALAREA 200.528 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 830.757 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNADIFFAREA 5.20755 LAYER metal4 ; 
    ANTENNAPARTIALMETALAREA 145.79 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 604.314 LAYER metal4 ;
  END DRAM_WEn[0]
  PIN DRAM_A[10] 
    ANTENNAPARTIALMETALAREA 122.43 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 507.21 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 90.5072 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 375.283 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.28045 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 77.896 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 323.037 LAYER metal5 ;
  END DRAM_A[10]
  PIN DRAM_A[9] 
    ANTENNAPARTIALMETALAREA 119.526 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 495.181 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 2.6656 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 11.368 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.25495 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 83.7648 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 347.35 LAYER metal5 ;
  END DRAM_A[9]
  PIN DRAM_A[8] 
    ANTENNAPARTIALMETALAREA 0.42 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.74 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 2.1616 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 9.28 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.25495 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 205.318 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 850.93 LAYER metal5 ;
  END DRAM_A[8]
  PIN DRAM_A[7] 
    ANTENNAPARTIALMETALAREA 7.3948 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 30.6356 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 31.1864 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 129.526 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.25495 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 197.994 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 820.584 LAYER metal5 ;
  END DRAM_A[7]
  PIN DRAM_A[6] 
    ANTENNAPARTIALMETALAREA 0.3976 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6472 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 2.0048 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 8.6304 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.25495 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 205.111 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 850.071 LAYER metal5 ;
  END DRAM_A[6]
  PIN DRAM_A[5] 
    ANTENNAPARTIALMETALAREA 0.3752 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.4368 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1344 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.25495 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 207.407 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 859.583 LAYER metal5 ;
  END DRAM_A[5]
  PIN DRAM_A[4] 
    ANTENNAPARTIALMETALAREA 0.4648 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9256 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 7.9632 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 33.3152 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.25495 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 200.67 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 831.674 LAYER metal5 ;
  END DRAM_A[4]
  PIN DRAM_A[3] 
    ANTENNAPARTIALMETALAREA 7.798 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 32.306 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 16.9176 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 70.412 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.25495 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 183.932 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 762.329 LAYER metal5 ;
  END DRAM_A[3]
  PIN DRAM_A[2] 
    ANTENNAPARTIALMETALAREA 3.2228 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.3516 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 47.32 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 196.365 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.25495 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 196.778 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 815.55 LAYER metal5 ;
  END DRAM_A[2]
  PIN DRAM_A[1] 
    ANTENNAPARTIALMETALAREA 2.6404 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.9388 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 55.3168 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 229.494 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.25495 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 209.104 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 866.613 LAYER metal5 ;
  END DRAM_A[1]
  PIN DRAM_A[0] 
    ANTENNAPARTIALMETALAREA 7.7756 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 32.2132 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 69.4456 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 288.028 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.25495 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 204.316 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 846.777 LAYER metal5 ;
  END DRAM_A[0]
  PIN DRAM_D[31] 
    ANTENNAPARTIALMETALAREA 7.3528 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 30.4616 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 74.3064 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 308.166 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 3.3804 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 192.752 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 798.869 LAYER metal5 ;
  END DRAM_D[31]
  PIN DRAM_D[30] 
    ANTENNAPARTIALMETALAREA 7.1092 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 29.4524 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 17.6848 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 73.5904 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.5386 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 180.841 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 749.522 LAYER metal5 ;
  END DRAM_D[30]
  PIN DRAM_D[29] 
    ANTENNAPARTIALMETALAREA 0.4732 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.9604 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 1.848 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 7.9808 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.5386 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 191.537 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 793.834 LAYER metal5 ;
  END DRAM_D[29]
  PIN DRAM_D[28] 
    ANTENNAPARTIALMETALAREA 0.4088 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.6936 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 3.1024 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 13.1776 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 3.3804 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 201.499 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 835.107 LAYER metal5 ;
  END DRAM_D[28]
  PIN DRAM_D[27] 
    ANTENNAPARTIALMETALAREA 0.5012 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0764 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1368 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.5386 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 194.208 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 804.901 LAYER metal5 ;
  END DRAM_D[27]
  PIN DRAM_D[26] 
    ANTENNAPARTIALMETALAREA 3.3516 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.8852 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 47.9472 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 198.963 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.5386 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 190.047 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 787.663 LAYER metal5 ;
  END DRAM_D[26]
  PIN DRAM_D[25] 
    ANTENNAPARTIALMETALAREA 2.5928 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.7416 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 71.4672 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 296.403 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 3.3804 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 187.718 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 778.012 LAYER metal5 ;
  END DRAM_D[25]
  PIN DRAM_D[24] 
    ANTENNAPARTIALMETALAREA 8.2348 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 34.1156 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 86.6936 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 359.484 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.5386 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 184.559 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 764.927 LAYER metal5 ;
  END DRAM_D[24]
  PIN DRAM_D[23] 
    ANTENNAPARTIALMETALAREA 7.6552 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 31.7144 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 106.904 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 443.213 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.6902 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 182.515 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 756.459 LAYER metal5 ;
  END DRAM_D[23]
  PIN DRAM_D[22] 
    ANTENNAPARTIALMETALAREA 8.0948 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 33.5356 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 128.106 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 531.048 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 3.3804 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 187.55 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 777.316 LAYER metal5 ;
  END DRAM_D[22]
  PIN DRAM_D[21] 
    ANTENNAPARTIALMETALAREA 7.336 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 30.392 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 156.8 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 649.925 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 3.3804 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 191.744 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 794.693 LAYER metal5 ;
  END DRAM_D[21]
  PIN DRAM_D[20] 
    ANTENNAPARTIALMETALAREA 0.364 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.508 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1368 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.6902 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 189.694 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 786.202 LAYER metal5 ;
  END DRAM_D[20]
  PIN DRAM_D[19] 
    ANTENNAPARTIALMETALAREA 6.3224 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 26.1928 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 205.061 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 849.862 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 3.3804 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 180.757 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 749.174 LAYER metal5 ;
  END DRAM_D[19]
  PIN DRAM_D[18] 
    ANTENNAPARTIALMETALAREA 5.5636 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 23.0492 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 219.957 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 911.574 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.6902 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 200.463 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 830.815 LAYER metal5 ;
  END DRAM_D[18]
  PIN DRAM_D[17] 
    ANTENNAPARTIALMETALAREA 4.9616 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 20.5552 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 235.323 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 975.235 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNADIFFAREA 1.6902 LAYER metal5 ; 
    ANTENNAPARTIALMETALAREA 185.618 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 769.312 LAYER metal5 ;
  END DRAM_D[17]
  PIN DRAM_D[16] 
    ANTENNAPARTIALMETALAREA 198.926 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 824.447 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNADIFFAREA 1.6902 LAYER metal4 ; 
    ANTENNAPARTIALMETALAREA 260.725 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1080.47 LAYER metal4 ;
  END DRAM_D[16]
  PIN DRAM_D[15] 
    ANTENNAPARTIALMETALAREA 0.5712 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3664 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNADIFFAREA 1.6902 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 1.8592 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.0272 LAYER metal3 ;
  END DRAM_D[15]
  PIN DRAM_D[14] 
    ANTENNAPARTIALMETALAREA 122.685 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 508.59 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNADIFFAREA 1.6902 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 53.732 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 222.929 LAYER metal3 ;
  END DRAM_D[14]
  PIN DRAM_D[13] 
    ANTENNADIFFAREA 1.6902 LAYER metal2 ; 
    ANTENNAPARTIALMETALAREA 409.245 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1696.09 LAYER metal2 ;
  END DRAM_D[13]
  PIN DRAM_D[12] 
    ANTENNADIFFAREA 1.6902 LAYER metal2 ; 
    ANTENNAPARTIALMETALAREA 402.889 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1669.76 LAYER metal2 ;
  END DRAM_D[12]
  PIN DRAM_D[11] 
    ANTENNAPARTIALMETALAREA 121.671 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 504.066 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNADIFFAREA 1.6902 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 109.11 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 452.354 LAYER metal3 ;
  END DRAM_D[11]
  PIN DRAM_D[10] 
    ANTENNADIFFAREA 1.5386 LAYER metal2 ; 
    ANTENNAPARTIALMETALAREA 400.302 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1659.04 LAYER metal2 ;
  END DRAM_D[10]
  PIN DRAM_D[9] 
    ANTENNADIFFAREA 1.5386 LAYER metal2 ; 
    ANTENNAPARTIALMETALAREA 397.39 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1646.98 LAYER metal2 ;
  END DRAM_D[9]
  PIN DRAM_D[8] 
    ANTENNADIFFAREA 1.5386 LAYER metal2 ; 
    ANTENNAPARTIALMETALAREA 397.351 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1646.82 LAYER metal2 ;
  END DRAM_D[8]
  PIN DRAM_D[7] 
    ANTENNAPARTIALMETALAREA 7.3212 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 30.218 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNADIFFAREA 1.6902 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 60.592 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 251.674 LAYER metal3 ;
  END DRAM_D[7]
  PIN DRAM_D[6] 
    ANTENNAPARTIALMETALAREA 7.3304 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 30.3688 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNADIFFAREA 1.6902 LAYER metal3 ; 
    ANTENNAPARTIALMETALAREA 7.9184 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 33.1296 LAYER metal3 ;
  END DRAM_D[6]
  PIN DRAM_D[5] 
    ANTENNADIFFAREA 3.3804 LAYER metal2 ; 
    ANTENNAPARTIALMETALAREA 397.298 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1646.27 LAYER metal2 ;
  END DRAM_D[5]
  PIN DRAM_D[4] 
    ANTENNADIFFAREA 3.3804 LAYER metal2 ; 
    ANTENNAPARTIALMETALAREA 398.294 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1650.08 LAYER metal2 ;
  END DRAM_D[4]
  PIN DRAM_D[3] 
    ANTENNADIFFAREA 1.5386 LAYER metal2 ; 
    ANTENNAPARTIALMETALAREA 181.563 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 752.19 LAYER metal2 ;
  END DRAM_D[3]
  PIN DRAM_D[2] 
    ANTENNADIFFAREA 1.5386 LAYER metal2 ; 
    ANTENNAPARTIALMETALAREA 181.048 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 750.381 LAYER metal2 ;
  END DRAM_D[2]
  PIN DRAM_D[1] 
    ANTENNADIFFAREA 1.5386 LAYER metal2 ; 
    ANTENNAPARTIALMETALAREA 208.225 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 862.97 LAYER metal2 ;
  END DRAM_D[1]
  PIN DRAM_D[0] 
    ANTENNADIFFAREA 1.5386 LAYER metal2 ; 
    ANTENNAPARTIALMETALAREA 398.311 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1650.8 LAYER metal2 ;
  END DRAM_D[0]
  PIN DRAM_Q[31] 
    ANTENNAPARTIALMETALAREA 0.3556 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4732 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 9.1504 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 38.2336 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 410.95 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1702.83 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.5936 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1088 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3186 LAYER metal5 ; 
    ANTENNAMAXAREACAR 367.647 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 1518.95 LAYER metal5 ;
    ANTENNAMAXCUTCAR 1.48205 LAYER via5 ;
  END DRAM_Q[31]
  PIN DRAM_Q[30] 
    ANTENNAPARTIALMETALAREA 2.6424 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.8344 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 68.1744 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 282.762 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4848 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1794.34 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5985.92 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3186 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5669.94 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18921 LAYER metal6 ;
  END DRAM_Q[30]
  PIN DRAM_Q[29] 
    ANTENNAPARTIALMETALAREA 3.2164 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 13.2124 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 52.8976 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 219.472 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4848 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1727.23 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5767.04 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3186 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5446.27 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18178.2 LAYER metal6 ;
  END DRAM_Q[29]
  PIN DRAM_Q[28] 
    ANTENNAPARTIALMETALAREA 7.1876 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 29.7772 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 29.9824 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 124.538 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.5936 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.784 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1717.63 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5730.24 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3186 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5430.72 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18140.6 LAYER metal6 ;
  END DRAM_Q[28]
  PIN DRAM_Q[27] 
    ANTENNAPARTIALMETALAREA 7.7392 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 32.0624 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 11.928 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 49.7408 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4848 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1705.06 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5693.12 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3186 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5400.26 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18066.1 LAYER metal6 ;
  END DRAM_Q[27]
  PIN DRAM_Q[26] 
    ANTENNAPARTIALMETALAREA 0.5712 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3664 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 1.8004 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.7836 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1368 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1729.15 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5768.64 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3186 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5476.31 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18309 LAYER metal6 ;
  END DRAM_Q[26]
  PIN DRAM_Q[25] 
    ANTENNAPARTIALMETALAREA 2.296 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.512 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 18.8776 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 78.532 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4848 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1733.86 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5784.32 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3186 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5456.51 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18202.6 LAYER metal6 ;
  END DRAM_Q[25]
  PIN DRAM_Q[24] 
    ANTENNAPARTIALMETALAREA 2.6704 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.9504 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 13.664 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 56.9328 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4848 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1721.09 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5741.76 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3186 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5441.15 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18174.1 LAYER metal6 ;
  END DRAM_Q[24]
  PIN DRAM_Q[23] 
    ANTENNAPARTIALMETALAREA 4.3344 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.9568 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.5712 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.6912 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4848 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1702.94 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5681.28 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3564 LAYER metal6 ; 
    ANTENNAMAXAREACAR 4829.41 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 16147.6 LAYER metal6 ;
  END DRAM_Q[23]
  PIN DRAM_Q[22] 
    ANTENNAPARTIALMETALAREA 4.3344 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.9568 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 8.302 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 34.7188 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4848 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1704.29 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5685.76 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3186 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5399.04 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18042.3 LAYER metal6 ;
  END DRAM_Q[22]
  PIN DRAM_Q[21] 
    ANTENNAPARTIALMETALAREA 4.3344 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.9568 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.6104 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.8536 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4848 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1700.26 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5672.32 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3186 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5365.04 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 17918.4 LAYER metal6 ;
  END DRAM_Q[21]
  PIN DRAM_Q[20] 
    ANTENNAPARTIALMETALAREA 5.9892 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 24.8124 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 1.3384 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.8696 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1368 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1725.02 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5754.88 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3186 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5437.35 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18153 LAYER metal6 ;
  END DRAM_Q[20]
  PIN DRAM_Q[19] 
    ANTENNAPARTIALMETALAREA 0.5712 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.3664 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.2632 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4152 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1368 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1368 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1741.92 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5811.2 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3186 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5495.24 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18328.7 LAYER metal6 ;
  END DRAM_Q[19]
  PIN DRAM_Q[18] 
    ANTENNAPARTIALMETALAREA 2.7664 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 11.4608 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 4.312 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 18.1888 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1368 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 1.6856 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 7.308 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1707.65 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5696.96 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3186 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5431.48 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18174.8 LAYER metal6 ;
  END DRAM_Q[18]
  PIN DRAM_Q[17] 
    ANTENNAPARTIALMETALAREA 7.3136 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 30.2992 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 12.0064 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 50.0656 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.4368 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1344 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1711.01 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5708.16 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3186 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5391.32 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 17997.9 LAYER metal6 ;
  END DRAM_Q[17]
  PIN DRAM_Q[16] 
    ANTENNAPARTIALMETALAREA 4.3288 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 17.9336 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 24.948 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 103.681 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.4368 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1344 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1728.1 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5765.12 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3186 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5464.85 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18252.4 LAYER metal6 ;
  END DRAM_Q[16]
  PIN DRAM_Q[15] 
    ANTENNAPARTIALMETALAREA 3.502 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 14.3956 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 48.0368 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 199.334 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4848 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1731.74 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5777.28 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3186 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5455.49 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18206.9 LAYER metal6 ;
  END DRAM_Q[15]
  PIN DRAM_Q[14] 
    ANTENNAPARTIALMETALAREA 4.8124 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 19.8244 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 72.3408 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 300.022 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4848 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1719.74 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5737.28 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3186 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5443.84 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18198.3 LAYER metal6 ;
  END DRAM_Q[14]
  PIN DRAM_Q[13] 
    ANTENNAPARTIALMETALAREA 3.836 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 15.892 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 88.6592 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 367.627 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4848 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.196 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.1368 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1722.29 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5755.36 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3186 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5465.98 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18307.1 LAYER metal6 ;
  END DRAM_Q[13]
  PIN DRAM_Q[12] 
    ANTENNAPARTIALMETALAREA 3.026 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.4236 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 124.594 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 516.502 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.4368 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.1344 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1730.5 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5773.12 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3186 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5459.39 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18223.7 LAYER metal6 ;
  END DRAM_Q[12]
  PIN DRAM_Q[11] 
    ANTENNAPARTIALMETALAREA 2.296 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.512 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 139.418 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 577.912 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4848 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1726.99 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5771.04 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3186 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5476.36 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18342.8 LAYER metal6 ;
  END DRAM_Q[11]
  PIN DRAM_Q[10] 
    ANTENNAPARTIALMETALAREA 7.9408 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 32.8976 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 38.7856 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 161.008 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4848 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1710.19 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5715.04 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3186 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5403 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18073.8 LAYER metal6 ;
  END DRAM_Q[10]
  PIN DRAM_Q[9] 
    ANTENNAPARTIALMETALAREA 7.6328 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 31.6216 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 173.863 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 720.615 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.5936 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.784 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1690.75 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5640.64 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3186 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5339.52 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 17829.5 LAYER metal6 ;
  END DRAM_Q[9]
  PIN DRAM_Q[8] 
    ANTENNAPARTIALMETALAREA 7.31 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 30.1716 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 192.125 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 796.27 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4848 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNADIFFAREA 0.36 LAYER metal6 ; 
    ANTENNAPARTIALMETALAREA 1719.5 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 5746.08 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3186 LAYER metal6 ; 
    ANTENNAMAXAREACAR 5441.85 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 18209.2 LAYER metal6 ;
  END DRAM_Q[8]
  PIN DRAM_Q[7] 
    ANTENNAPARTIALMETALAREA 2.6004 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.6604 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 14.532 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 60.5288 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 393.081 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1628.8 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.5936 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1088 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3186 LAYER metal5 ; 
    ANTENNAMAXAREACAR 42.7868 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 166.81 LAYER metal5 ;
    ANTENNAMAXCUTCAR 1.23318 LAYER via5 ;
  END DRAM_Q[7]
  PIN DRAM_Q[6] 
    ANTENNAPARTIALMETALAREA 2.296 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.512 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 0.8904 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.6632 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 4.3568 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 18.3744 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3564 LAYER metal4 ; 
    ANTENNAMAXAREACAR 34.7299 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 130.545 LAYER metal4 ;
    ANTENNAMAXCUTCAR 0.934905 LAYER via4 ;
  END DRAM_Q[6]
  PIN DRAM_Q[5] 
    ANTENNAPARTIALMETALAREA 6.7172 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 28.1532 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 64.7752 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 268.679 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 299.69 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1241.9 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNAPARTIALMETALAREA 18 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 69.6 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3564 LAYER metal6 ; 
    ANTENNAMAXAREACAR 108.914 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 430.31 LAYER metal6 ;
  END DRAM_Q[5]
  PIN DRAM_Q[4] 
    ANTENNAPARTIALMETALAREA 3.0996 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.166 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 21.448 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 89.1808 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 282.072 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1168.91 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNAPARTIALMETALAREA 18 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 69.6 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3564 LAYER metal6 ; 
    ANTENNAMAXAREACAR 89.0652 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 352.108 LAYER metal6 ;
  END DRAM_Q[4]
  PIN DRAM_Q[3] 
    ANTENNAPARTIALMETALAREA 6.7956 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 28.1532 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 353.427 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1464.52 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 4.8496 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 21.0656 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3186 LAYER metal5 ; 
    ANTENNAMAXAREACAR 75.4155 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 310.31 LAYER metal5 ;
    ANTENNAMAXCUTCAR 1.96032 LAYER via5 ;
  END DRAM_Q[3]
  PIN DRAM_Q[2] 
    ANTENNAPARTIALMETALAREA 6.0956 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 25.2532 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 336.65 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1395.34 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.5936 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1088 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3564 LAYER metal5 ; 
    ANTENNAMAXAREACAR 34.2036 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 130.415 LAYER metal5 ;
    ANTENNAMAXCUTCAR 1.42985 LAYER via5 ;
  END DRAM_Q[2]
  PIN DRAM_Q[1] 
    ANTENNAPARTIALMETALAREA 4.2784 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.024 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3564 LAYER metal3 ; 
    ANTENNAMAXAREACAR 42.658 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 175.439 LAYER metal3 ;
    ANTENNAMAXCUTCAR 1.18788 LAYER via3 ;
  END DRAM_Q[1]
  PIN DRAM_Q[0] 
    ANTENNAPARTIALMETALAREA 7.6412 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 31.6564 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 292.242 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1211.36 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.5936 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1088 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3186 LAYER metal5 ; 
    ANTENNAMAXAREACAR 25.1222 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 92.3188 LAYER metal5 ;
    ANTENNAMAXCUTCAR 1.48205 LAYER via5 ;
  END DRAM_Q[0]
  PIN sensor_out[31] 
    ANTENNAPARTIALMETALAREA 2.1252 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.454 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1962 LAYER metal3 ; 
    ANTENNAMAXAREACAR 33.5882 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 138.135 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.799185 LAYER via3 ;
  END sensor_out[31]
  PIN sensor_out[30] 
    ANTENNAPARTIALMETALAREA 1.1956 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.9276 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1584 LAYER metal3 ; 
    ANTENNAMAXAREACAR 40.6831 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 161.816 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.989899 LAYER via3 ;
  END sensor_out[30]
  PIN sensor_out[29] 
    ANTENNAPARTIALMETALAREA 4.144 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 18.1424 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1584 LAYER metal3 ; 
    ANTENNAMAXAREACAR 50.6705 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 201.141 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.989899 LAYER via3 ;
  END sensor_out[29]
  PIN sensor_out[28] 
    ANTENNAPARTIALMETALAREA 0.3668 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5196 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 162.568 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 674.146 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.5936 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1088 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4188 LAYER metal5 ; 
    ANTENNAMAXAREACAR 10.9637 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 45.3257 LAYER metal5 ;
    ANTENNAMAXCUTCAR 0.748806 LAYER via5 ;
  END sensor_out[28]
  PIN sensor_out[27] 
    ANTENNAPARTIALMETALAREA 1.022 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.234 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 131.992 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 547.149 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.5936 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1088 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4188 LAYER metal5 ; 
    ANTENNAMAXAREACAR 16.1385 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 69.0907 LAYER metal5 ;
    ANTENNAMAXCUTCAR 0.748806 LAYER via5 ;
  END sensor_out[27]
  PIN sensor_out[26] 
    ANTENNAPARTIALMETALAREA 348.723 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1445.04 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 2.7888 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 11.8784 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4188 LAYER metal4 ; 
    ANTENNAMAXAREACAR 9.84814 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 39.0067 LAYER metal4 ;
    ANTENNAMAXCUTCAR 0.561605 LAYER via4 ;
  END sensor_out[26]
  PIN sensor_out[25] 
    ANTENNAPARTIALMETALAREA 170.713 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 707.565 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 4.3232 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 18.8848 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1584 LAYER metal4 ; 
    ANTENNAMAXAREACAR 36.423 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 144.167 LAYER metal4 ;
    ANTENNAMAXCUTCAR 1.48485 LAYER via4 ;
  END sensor_out[25]
  PIN sensor_out[24] 
    ANTENNAPARTIALMETALAREA 5.306 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 22.3068 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 2.4752 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 10.5792 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.5936 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1088 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1584 LAYER metal5 ; 
    ANTENNAMAXAREACAR 40.2058 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 163.939 LAYER metal5 ;
    ANTENNAMAXCUTCAR 1.9798 LAYER via5 ;
  END sensor_out[24]
  PIN sensor_out[23] 
    ANTENNAPARTIALMETALAREA 178.872 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 741.368 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.56 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9696 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1584 LAYER metal4 ; 
    ANTENNAMAXAREACAR 38.9331 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 152.515 LAYER metal4 ;
    ANTENNAMAXCUTCAR 1.48485 LAYER via4 ;
  END sensor_out[23]
  PIN sensor_out[22] 
    ANTENNAPARTIALMETALAREA 13.3896 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 56.1208 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1584 LAYER metal3 ; 
    ANTENNAMAXAREACAR 93.7664 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 377.631 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.989899 LAYER via3 ;
  END sensor_out[22]
  PIN sensor_out[21] 
    ANTENNAPARTIALMETALAREA 0.8428 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.4916 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1584 LAYER metal3 ; 
    ANTENNAMAXAREACAR 79.2348 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 322.21 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.989899 LAYER via3 ;
  END sensor_out[21]
  PIN sensor_out[20] 
    ANTENNAPARTIALMETALAREA 78.4364 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 324.951 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal3 ; 
    ANTENNAMAXAREACAR 253.981 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 1047.21 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.500639 LAYER via3 ;
  END sensor_out[20]
  PIN sensor_out[19] 
    ANTENNAPARTIALMETALAREA 11.8552 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 49.4392 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal3 ; 
    ANTENNAMAXAREACAR 58.8129 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 240.733 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.500639 LAYER via3 ;
  END sensor_out[19]
  PIN sensor_out[18] 
    ANTENNAPARTIALMETALAREA 149.248 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 618.64 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.56 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9696 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1584 LAYER metal4 ; 
    ANTENNAMAXAREACAR 17.6149 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 64.197 LAYER metal4 ;
    ANTENNAMAXCUTCAR 1.48485 LAYER via4 ;
  END sensor_out[18]
  PIN sensor_out[17] 
    ANTENNAPARTIALMETALAREA 156.825 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 650.029 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 4.2336 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 17.864 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1584 LAYER metal4 ; 
    ANTENNAMAXAREACAR 38.1907 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 147.389 LAYER metal4 ;
    ANTENNAMAXCUTCAR 1.48485 LAYER via4 ;
  END sensor_out[17]
  PIN sensor_out[16] 
    ANTENNAPARTIALMETALAREA 3.6064 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.9408 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal3 ; 
    ANTENNAMAXAREACAR 118.693 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 487.77 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.500639 LAYER via3 ;
  END sensor_out[16]
  PIN sensor_out[15] 
    ANTENNAPARTIALMETALAREA 0.6636 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.7492 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 1.6912 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 7.3312 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.5936 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 3.1088 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4188 LAYER metal5 ; 
    ANTENNAMAXAREACAR 391.468 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 1623.01 LAYER metal5 ;
    ANTENNAMAXCUTCAR 0.748806 LAYER via5 ;
  END sensor_out[15]
  PIN sensor_out[14] 
    ANTENNAPARTIALMETALAREA 154.535 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 640.54 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4848 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 4.9672 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 20.9032 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1584 LAYER metal5 ; 
    ANTENNAMAXAREACAR 55.4432 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 220.914 LAYER metal5 ;
    ANTENNAMAXCUTCAR 1.9798 LAYER via5 ;
  END sensor_out[14]
  PIN sensor_out[13] 
    ANTENNAPARTIALMETALAREA 158.925 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 658.729 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4188 LAYER metal3 ; 
    ANTENNAMAXAREACAR 391.939 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 1621.32 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.374403 LAYER via3 ;
  END sensor_out[13]
  PIN sensor_out[12] 
    ANTENNAPARTIALMETALAREA 149.377 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 619.173 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.56 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 2.9696 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1584 LAYER metal4 ; 
    ANTENNAMAXAREACAR 17.0492 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 61.8535 LAYER metal4 ;
    ANTENNAMAXCUTCAR 1.48485 LAYER via4 ;
  END sensor_out[12]
  PIN sensor_out[11] 
    ANTENNAPARTIALMETALAREA 156.965 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 650.609 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4848 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 4.2896 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 18.096 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1584 LAYER metal5 ; 
    ANTENNAMAXAREACAR 70.6099 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 283.747 LAYER metal5 ;
    ANTENNAMAXCUTCAR 1.9798 LAYER via5 ;
  END sensor_out[11]
  PIN sensor_out[10] 
    ANTENNAPARTIALMETALAREA 157.349 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 652.198 LAYER metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4188 LAYER metal3 ; 
    ANTENNAMAXAREACAR 391.13 LAYER metal3 ;
    ANTENNAMAXSIDEAREACAR 1617.97 LAYER metal3 ;
    ANTENNAMAXCUTCAR 0.374403 LAYER via3 ;
  END sensor_out[10]
  PIN sensor_out[9] 
    ANTENNAPARTIALMETALAREA 5.278 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 22.1908 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 7.1792 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 30.0672 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 5.544 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 23.9424 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1584 LAYER metal5 ; 
    ANTENNAMAXAREACAR 64.8472 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 266.025 LAYER metal5 ;
    ANTENNAMAXCUTCAR 1.9798 LAYER via5 ;
  END sensor_out[9]
  PIN sensor_out[8] 
    ANTENNAPARTIALMETALAREA 151.312 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 627.189 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 0.28 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.4848 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 4.9504 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 20.8336 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1584 LAYER metal5 ; 
    ANTENNAMAXAREACAR 70.2765 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 284.03 LAYER metal5 ;
    ANTENNAMAXCUTCAR 1.9798 LAYER via5 ;
  END sensor_out[8]
  PIN sensor_out[7] 
    ANTENNAPARTIALMETALAREA 6.4148 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 26.5756 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 217.134 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 899.882 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 321.91 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1333.95 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNAPARTIALMETALAREA 53.184 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 182.08 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4188 LAYER metal6 ; 
    ANTENNAMAXAREACAR 137.18 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 476.103 LAYER metal6 ;
  END sensor_out[7]
  PIN sensor_out[6] 
    ANTENNAPARTIALMETALAREA 7.8092 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 32.3524 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 235.95 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 977.834 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 288.266 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1194.57 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNAPARTIALMETALAREA 62.592 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 213.44 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4188 LAYER metal6 ; 
    ANTENNAMAXAREACAR 157.63 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 542.3 LAYER metal6 ;
  END sensor_out[6]
  PIN sensor_out[5] 
    ANTENNAPARTIALMETALAREA 6.9412 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 28.7564 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 264.331 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1095.41 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 287.414 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1191.04 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNAPARTIALMETALAREA 23.616 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 83.52 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4188 LAYER metal6 ; 
    ANTENNAMAXAREACAR 101.946 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 388.063 LAYER metal6 ;
  END sensor_out[5]
  PIN sensor_out[4] 
    ANTENNAPARTIALMETALAREA 5.9108 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 24.4876 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 297.259 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1231.83 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 297.276 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1231.9 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNAPARTIALMETALAREA 18 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 69.6 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4188 LAYER metal6 ; 
    ANTENNAMAXAREACAR 52.3391 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 204.092 LAYER metal6 ;
  END sensor_out[4]
  PIN sensor_out[3] 
    ANTENNAPARTIALMETALAREA 1.75 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.25 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 306.981 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1272.1 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNAPARTIALMETALAREA 17.568 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 63.36 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4188 LAYER metal6 ; 
    ANTENNAMAXAREACAR 58.4613 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 221.931 LAYER metal6 ;
  END sensor_out[3]
  PIN sensor_out[2] 
    ANTENNAPARTIALMETALAREA 6.79 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 28.13 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 327.712 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1357.99 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 290.382 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1203.34 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNAPARTIALMETALAREA 51.168 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 175.36 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4188 LAYER metal6 ; 
    ANTENNAMAXAREACAR 126.255 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 434.741 LAYER metal6 ;
  END sensor_out[2]
  PIN sensor_out[1] 
    ANTENNAPARTIALMETALAREA 7.49 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 31.03 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 348.88 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1445.68 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 316.389 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1311.08 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNAPARTIALMETALAREA 58.56 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 200 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4188 LAYER metal6 ; 
    ANTENNAMAXAREACAR 146.887 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 505.929 LAYER metal6 ;
  END sensor_out[1]
  PIN sensor_out[0] 
    ANTENNAPARTIALMETALAREA 1.386 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.742 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 373.688 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1548.46 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNAPARTIALMETALAREA 17.568 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 63.36 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.068 LAYER metal6 ; 
    ANTENNAMAXAREACAR 27.3635 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 103.541 LAYER metal6 ;
  END sensor_out[0]
  PIN clk 
    ANTENNAPARTIALMETALAREA 0.728 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.016 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 133.448 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 553.181 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 217.448 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 901.181 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.3622 LAYER metal4 ; 
    ANTENNAMAXAREACAR 41.895 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 168.656 LAYER metal4 ;
    ANTENNAMAXCUTCAR 0.0438626 LAYER via4 ;
  END clk
  PIN clk2 
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 78.344 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 324.893 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 220.898 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 915.472 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 5.3622 LAYER metal4 ; 
    ANTENNAMAXAREACAR 42.5384 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 171.321 LAYER metal4 ;
    ANTENNAMAXCUTCAR 0.0438626 LAYER via4 ;
  END clk2
  PIN rst 
    ANTENNAPARTIALMETALAREA 1.9824 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 8.2128 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 36.12 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 149.965 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 25.6984 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 106.79 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3132 LAYER metal4 ; 
    ANTENNAMAXAREACAR 86.8844 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 357.029 LAYER metal4 ;
    ANTENNAMAXCUTCAR 0.750958 LAYER via4 ;
  END rst
  PIN rst2 
    ANTENNAPARTIALMETALAREA 7.3136 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 30.2992 LAYER metal2 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via2 ;
    ANTENNAPARTIALMETALAREA 193.346 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 801.328 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 389.463 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1613.82 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 0.2968 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.5544 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNAPARTIALMETALAREA 20.256 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 72.32 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1962 LAYER metal6 ; 
    ANTENNAMAXAREACAR 119.89 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 439.87 LAYER metal6 ;
  END rst2
  PIN DRAM_valid 
    ANTENNAPARTIALMETALAREA 7.1204 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 29.4988 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 262.293 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1086.97 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 5.2304 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 22.6432 LAYER metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.2642 LAYER metal5 ; 
    ANTENNAMAXAREACAR 229.094 LAYER metal5 ;
    ANTENNAMAXSIDEAREACAR 947.658 LAYER metal5 ;
    ANTENNAMAXCUTCAR 2.79715 LAYER via5 ;
  END DRAM_valid
  PIN sensor_ready 
    ANTENNAPARTIALMETALAREA 7.9772 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 33.0484 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNAPARTIALMETALAREA 249.312 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1033.19 LAYER metal4 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via4 ;
    ANTENNAPARTIALMETALAREA 325.416 LAYER metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1348.48 LAYER metal5 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via5 ;
    ANTENNAPARTIALMETALAREA 18 LAYER metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 69.6 LAYER metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1584 LAYER metal6 ; 
    ANTENNAMAXAREACAR 162.343 LAYER metal6 ;
    ANTENNAMAXSIDEAREACAR 641.283 LAYER metal6 ;
  END sensor_ready
  PIN ROM_enable 
    ANTENNADIFFAREA 1.5386 LAYER metal2 ; 
    ANTENNAPARTIALMETALAREA 122.296 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 507.303 LAYER metal2 ;
  END ROM_enable
  PIN ROM_read 
    ANTENNADIFFAREA 1.5386 LAYER metal2 ; 
    ANTENNAPARTIALMETALAREA 142.019 LAYER metal2 ;
    ANTENNAPARTIALMETALSIDEAREA 589.013 LAYER metal2 ;
  END ROM_read
  PIN DRAM_CSn 
    ANTENNAPARTIALMETALAREA 209.868 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 869.455 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNADIFFAREA 1.0927 LAYER metal4 ; 
    ANTENNAPARTIALMETALAREA 244.782 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1014.42 LAYER metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9708 LAYER metal4 ; 
    ANTENNAMAXAREACAR 263.703 LAYER metal4 ;
    ANTENNAMAXSIDEAREACAR 1088.49 LAYER metal4 ;
    ANTENNAMAXCUTCAR 0.748092 LAYER via4 ;
  END DRAM_CSn
  PIN DRAM_RASn 
    ANTENNAPARTIALMETALAREA 190.226 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 788.081 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNADIFFAREA 1.66835 LAYER metal4 ; 
    ANTENNAPARTIALMETALAREA 119.605 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 495.83 LAYER metal4 ;
  END DRAM_RASn
  PIN DRAM_CASn 
    ANTENNAPARTIALMETALAREA 199.284 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 825.607 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNADIFFAREA 1.66835 LAYER metal4 ; 
    ANTENNAPARTIALMETALAREA 105.666 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 438.086 LAYER metal4 ;
  END DRAM_CASn
  PIN sensor_en 
    ANTENNAPARTIALMETALAREA 0.42 LAYER metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.74 LAYER metal3 ;
    ANTENNAPARTIALCUTAREA 0.0784 LAYER via3 ;
    ANTENNADIFFAREA 1.5386 LAYER metal4 ; 
    ANTENNAPARTIALMETALAREA 404.387 LAYER metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1675.64 LAYER metal4 ;
  END sensor_en
END top

END LIBRARY
